** Profile: "SCHEMATIC1-Task_1"  [ C:\Users\Asad Ur Rehman\Desktop\DC_DC_Converters\Task_1\Task_1-PSpiceFiles\SCHEMATIC1\Task_1.sim ] 

** Creating circuit file "Task_1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Asad Ur Rehman\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "C:\Users\Asad Ur Rehman\Desktop\ELEC4170_Fall_2024.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40m 0 1e-6 SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
